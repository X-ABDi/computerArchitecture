module alu (
    input [31:0] pc,
    input [31:0] 
);

endmodule